module multiplier(input [3:0] a, input [3:0] b, output [7:0] prod);
  assign prod = a * b;
endmodule
