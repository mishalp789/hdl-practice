module multiplier(input [3:0] a, b, output [7:0] product);
  assign product = a * b;
endmodule

