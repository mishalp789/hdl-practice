// Day 1: Hello World in SystemVerilog
